module Signal_ROM_2 (
    input clk,  // clock
    //input rst,  // reset
    output [7:0] Signal_out
  );
  localparam SIZE_b = 7'b1111110;//7'b1111110 <========= update here
  reg [7:0] signal_q;
  assign Signal_out = signal_q;
  reg [7:0]addr;
  reg [6:0] busy_counter = 7'b0;//7 bits
  reg [7:0] Signal [0:2][0:255];
  /*
assign Signal[0][0] = 8'b01001011; assign Signal[1][0] = 8'b00001011; assign Signal[2][0] = 8'b00011001; 
assign Signal[0][1] = 8'b01001100; assign Signal[1][1] = 8'b00001011; assign Signal[2][1] = 8'b00011001; 
assign Signal[0][2] = 8'b01001101; assign Signal[1][2] = 8'b00001100; assign Signal[2][2] = 8'b00011001; 
assign Signal[0][3] = 8'b01001110; assign Signal[1][3] = 8'b00001100; assign Signal[2][3] = 8'b00011001; 
assign Signal[0][4] = 8'b01001111; assign Signal[1][4] = 8'b00001100; assign Signal[2][4] = 8'b00011001; 
assign Signal[0][5] = 8'b01010001; assign Signal[1][5] = 8'b00001100; assign Signal[2][5] = 8'b00011001; 
assign Signal[0][6] = 8'b01010010; assign Signal[1][6] = 8'b00001100; assign Signal[2][6] = 8'b00011001; 
assign Signal[0][7] = 8'b01010011; assign Signal[1][7] = 8'b00001100; assign Signal[2][7] = 8'b00011001; 
assign Signal[0][8] = 8'b01010100; assign Signal[1][8] = 8'b00001100; assign Signal[2][8] = 8'b00011001; 
assign Signal[0][9] = 8'b01010101; assign Signal[1][9] = 8'b00001100; assign Signal[2][9] = 8'b00011001; 
assign Signal[0][10] = 8'b01010111; assign Signal[1][10] = 8'b00001101; assign Signal[2][10] = 8'b00011001; 
assign Signal[0][11] = 8'b01011000; assign Signal[1][11] = 8'b00001101; assign Signal[2][11] = 8'b00011001; 
assign Signal[0][12] = 8'b01011001; assign Signal[1][12] = 8'b00001101; assign Signal[2][12] = 8'b00011001; 
assign Signal[0][13] = 8'b01011010; assign Signal[1][13] = 8'b00001101; assign Signal[2][13] = 8'b00011001; 
assign Signal[0][14] = 8'b01011011; assign Signal[1][14] = 8'b00001101; assign Signal[2][14] = 8'b00011001; 
assign Signal[0][15] = 8'b01011100; assign Signal[1][15] = 8'b00001101; assign Signal[2][15] = 8'b00011001; 
assign Signal[0][16] = 8'b01011110; assign Signal[1][16] = 8'b00001101; assign Signal[2][16] = 8'b00011001; 
assign Signal[0][17] = 8'b01011111; assign Signal[1][17] = 8'b00001110; assign Signal[2][17] = 8'b00011001; 
assign Signal[0][18] = 8'b01100000; assign Signal[1][18] = 8'b00001110; assign Signal[2][18] = 8'b00011001; 
assign Signal[0][19] = 8'b01100001; assign Signal[1][19] = 8'b00001110; assign Signal[2][19] = 8'b00011001; 
assign Signal[0][20] = 8'b01100010; assign Signal[1][20] = 8'b00001110; assign Signal[2][20] = 8'b00011001; 
assign Signal[0][21] = 8'b01100011; assign Signal[1][21] = 8'b00001110; assign Signal[2][21] = 8'b00011001; 
assign Signal[0][22] = 8'b01100100; assign Signal[1][22] = 8'b00001110; assign Signal[2][22] = 8'b00011001; 
assign Signal[0][23] = 8'b01100101; assign Signal[1][23] = 8'b00001110; assign Signal[2][23] = 8'b00011001; 
assign Signal[0][24] = 8'b01100110; assign Signal[1][24] = 8'b00001111; assign Signal[2][24] = 8'b00011001; 
assign Signal[0][25] = 8'b01100111; assign Signal[1][25] = 8'b00001111; assign Signal[2][25] = 8'b00011001; 
assign Signal[0][26] = 8'b01101000; assign Signal[1][26] = 8'b00001111; assign Signal[2][26] = 8'b00011001; 
assign Signal[0][27] = 8'b01101001; assign Signal[1][27] = 8'b00001111; assign Signal[2][27] = 8'b00011001; 
assign Signal[0][28] = 8'b01101010; assign Signal[1][28] = 8'b00001111; assign Signal[2][28] = 8'b00011001; 
assign Signal[0][29] = 8'b01101011; assign Signal[1][29] = 8'b00001111; assign Signal[2][29] = 8'b00011001; 
assign Signal[0][30] = 8'b01101100; assign Signal[1][30] = 8'b00010000; assign Signal[2][30] = 8'b00011001; 
assign Signal[0][31] = 8'b01101101; assign Signal[1][31] = 8'b00010000; assign Signal[2][31] = 8'b00011001; 
assign Signal[0][32] = 8'b01101110; assign Signal[1][32] = 8'b00010000; assign Signal[2][32] = 8'b00011001; 
assign Signal[0][33] = 8'b01101111; assign Signal[1][33] = 8'b00010000; assign Signal[2][33] = 8'b00011001; 
assign Signal[0][34] = 8'b01110000; assign Signal[1][34] = 8'b00010000; assign Signal[2][34] = 8'b00011001; 
assign Signal[0][35] = 8'b01110000; assign Signal[1][35] = 8'b00010001; assign Signal[2][35] = 8'b00011010; 
assign Signal[0][36] = 8'b01110001; assign Signal[1][36] = 8'b00010001; assign Signal[2][36] = 8'b00011010; 
assign Signal[0][37] = 8'b01110010; assign Signal[1][37] = 8'b00010001; assign Signal[2][37] = 8'b00011010; 
assign Signal[0][38] = 8'b01110011; assign Signal[1][38] = 8'b00010001; assign Signal[2][38] = 8'b00011010; 
assign Signal[0][39] = 8'b01110011; assign Signal[1][39] = 8'b00010001; assign Signal[2][39] = 8'b00011010; 
assign Signal[0][40] = 8'b01110100; assign Signal[1][40] = 8'b00010010; assign Signal[2][40] = 8'b00011010; 
assign Signal[0][41] = 8'b01110101; assign Signal[1][41] = 8'b00010010; assign Signal[2][41] = 8'b00011010; 
assign Signal[0][42] = 8'b01110101; assign Signal[1][42] = 8'b00010010; assign Signal[2][42] = 8'b00011010; 
assign Signal[0][43] = 8'b01110110; assign Signal[1][43] = 8'b00010010; assign Signal[2][43] = 8'b00011010; 
assign Signal[0][44] = 8'b01110111; assign Signal[1][44] = 8'b00010011; assign Signal[2][44] = 8'b00011010; 
assign Signal[0][45] = 8'b01110111; assign Signal[1][45] = 8'b00010011; assign Signal[2][45] = 8'b00011010; 
assign Signal[0][46] = 8'b01111000; assign Signal[1][46] = 8'b00010011; assign Signal[2][46] = 8'b00011010; 
assign Signal[0][47] = 8'b01111000; assign Signal[1][47] = 8'b00010011; assign Signal[2][47] = 8'b00011010; 
assign Signal[0][48] = 8'b01111001; assign Signal[1][48] = 8'b00010100; assign Signal[2][48] = 8'b00011010; 
assign Signal[0][49] = 8'b01111001; assign Signal[1][49] = 8'b00010100; assign Signal[2][49] = 8'b00011011; 
assign Signal[0][50] = 8'b01111010; assign Signal[1][50] = 8'b00010100; assign Signal[2][50] = 8'b00011011; 
assign Signal[0][51] = 8'b01111010; assign Signal[1][51] = 8'b00010100; assign Signal[2][51] = 8'b00011011; 
assign Signal[0][52] = 8'b01111010; assign Signal[1][52] = 8'b00010101; assign Signal[2][52] = 8'b00011011; 
assign Signal[0][53] = 8'b01111011; assign Signal[1][53] = 8'b00010101; assign Signal[2][53] = 8'b00011011; 
assign Signal[0][54] = 8'b01111011; assign Signal[1][54] = 8'b00010101; assign Signal[2][54] = 8'b00011011; 
assign Signal[0][55] = 8'b01111011; assign Signal[1][55] = 8'b00010101; assign Signal[2][55] = 8'b00011011; 
assign Signal[0][56] = 8'b01111100; assign Signal[1][56] = 8'b00010110; assign Signal[2][56] = 8'b00011011; 
assign Signal[0][57] = 8'b01111100; assign Signal[1][57] = 8'b00010110; assign Signal[2][57] = 8'b00011011; 
assign Signal[0][58] = 8'b01111100; assign Signal[1][58] = 8'b00010110; assign Signal[2][58] = 8'b00011100; 
assign Signal[0][59] = 8'b01111100; assign Signal[1][59] = 8'b00010111; assign Signal[2][59] = 8'b00011100; 
assign Signal[0][60] = 8'b01111100; assign Signal[1][60] = 8'b00010111; assign Signal[2][60] = 8'b00011100; 
assign Signal[0][61] = 8'b01111100; assign Signal[1][61] = 8'b00010111; assign Signal[2][61] = 8'b00011100; 
assign Signal[0][62] = 8'b01111100; assign Signal[1][62] = 8'b00011000; assign Signal[2][62] = 8'b00011100; 
assign Signal[0][63] = 8'b01111100; assign Signal[1][63] = 8'b00011000; assign Signal[2][63] = 8'b00011100; 
assign Signal[0][64] = 8'b01111101; assign Signal[1][64] = 8'b00011000; assign Signal[2][64] = 8'b00011101; 
assign Signal[0][65] = 8'b01111100; assign Signal[1][65] = 8'b00011001; assign Signal[2][65] = 8'b00011101; 
assign Signal[0][66] = 8'b01111100; assign Signal[1][66] = 8'b00011001; assign Signal[2][66] = 8'b00011101; 
assign Signal[0][67] = 8'b01111100; assign Signal[1][67] = 8'b00011001; assign Signal[2][67] = 8'b00011101; 
assign Signal[0][68] = 8'b01111100; assign Signal[1][68] = 8'b00011010; assign Signal[2][68] = 8'b00011101; 
assign Signal[0][69] = 8'b01111100; assign Signal[1][69] = 8'b00011010; assign Signal[2][69] = 8'b00011110; 
assign Signal[0][70] = 8'b01111100; assign Signal[1][70] = 8'b00011011; assign Signal[2][70] = 8'b00011110; 
assign Signal[0][71] = 8'b01111100; assign Signal[1][71] = 8'b00011011; assign Signal[2][71] = 8'b00011110; 
assign Signal[0][72] = 8'b01111100; assign Signal[1][72] = 8'b00011011; assign Signal[2][72] = 8'b00011111; 
assign Signal[0][73] = 8'b01111011; assign Signal[1][73] = 8'b00011100; assign Signal[2][73] = 8'b00011111; 
assign Signal[0][74] = 8'b01111011; assign Signal[1][74] = 8'b00011100; assign Signal[2][74] = 8'b00011111; 
assign Signal[0][75] = 8'b01111011; assign Signal[1][75] = 8'b00011101; assign Signal[2][75] = 8'b00011111; 
assign Signal[0][76] = 8'b01111010; assign Signal[1][76] = 8'b00011101; assign Signal[2][76] = 8'b00100000; 
assign Signal[0][77] = 8'b01111010; assign Signal[1][77] = 8'b00011110; assign Signal[2][77] = 8'b00100000; 
assign Signal[0][78] = 8'b01111010; assign Signal[1][78] = 8'b00011110; assign Signal[2][78] = 8'b00100000; 
assign Signal[0][79] = 8'b01111001; assign Signal[1][79] = 8'b00011111; assign Signal[2][79] = 8'b00100001; 
assign Signal[0][80] = 8'b01111001; assign Signal[1][80] = 8'b00011111; assign Signal[2][80] = 8'b00100001; 
assign Signal[0][81] = 8'b01111000; assign Signal[1][81] = 8'b00100000; assign Signal[2][81] = 8'b00100010; 
assign Signal[0][82] = 8'b01111000; assign Signal[1][82] = 8'b00100000; assign Signal[2][82] = 8'b00100010; 
assign Signal[0][83] = 8'b01110111; assign Signal[1][83] = 8'b00100001; assign Signal[2][83] = 8'b00100010; 
assign Signal[0][84] = 8'b01110111; assign Signal[1][84] = 8'b00100001; assign Signal[2][84] = 8'b00100011; 
assign Signal[0][85] = 8'b01110110; assign Signal[1][85] = 8'b00100010; assign Signal[2][85] = 8'b00100011; 
assign Signal[0][86] = 8'b01110101; assign Signal[1][86] = 8'b00100010; assign Signal[2][86] = 8'b00100100; 
assign Signal[0][87] = 8'b01110101; assign Signal[1][87] = 8'b00100011; assign Signal[2][87] = 8'b00100100; 
assign Signal[0][88] = 8'b01110100; assign Signal[1][88] = 8'b00100100; assign Signal[2][88] = 8'b00100101; 
assign Signal[0][89] = 8'b01110011; assign Signal[1][89] = 8'b00100100; assign Signal[2][89] = 8'b00100101; 
assign Signal[0][90] = 8'b01110011; assign Signal[1][90] = 8'b00100101; assign Signal[2][90] = 8'b00100110; 
assign Signal[0][91] = 8'b01110010; assign Signal[1][91] = 8'b00100110; assign Signal[2][91] = 8'b00100110; 
assign Signal[0][92] = 8'b01110001; assign Signal[1][92] = 8'b00100110; assign Signal[2][92] = 8'b00100111; 
assign Signal[0][93] = 8'b01110000; assign Signal[1][93] = 8'b00100111; assign Signal[2][93] = 8'b00101000; 
assign Signal[0][94] = 8'b01110000; assign Signal[1][94] = 8'b00101000; assign Signal[2][94] = 8'b00101000; 
assign Signal[0][95] = 8'b01101111; assign Signal[1][95] = 8'b00101000; assign Signal[2][95] = 8'b00101001; 
assign Signal[0][96] = 8'b01101110; assign Signal[1][96] = 8'b00101001; assign Signal[2][96] = 8'b00101010; 
assign Signal[0][97] = 8'b01101101; assign Signal[1][97] = 8'b00101010; assign Signal[2][97] = 8'b00101010; 
assign Signal[0][98] = 8'b01101100; assign Signal[1][98] = 8'b00101011; assign Signal[2][98] = 8'b00101011; 
assign Signal[0][99] = 8'b01101011; assign Signal[1][99] = 8'b00101100; assign Signal[2][99] = 8'b00101100; 
assign Signal[0][100] = 8'b01101010; assign Signal[1][100] = 8'b00101100; assign Signal[2][100] = 8'b00101101; 
assign Signal[0][101] = 8'b01101001; assign Signal[1][101] = 8'b00101101; assign Signal[2][101] = 8'b00101101; 
assign Signal[0][102] = 8'b01101000; assign Signal[1][102] = 8'b00101110; assign Signal[2][102] = 8'b00101110; 
assign Signal[0][103] = 8'b01100111; assign Signal[1][103] = 8'b00101111; assign Signal[2][103] = 8'b00101111; 
assign Signal[0][104] = 8'b01100110; assign Signal[1][104] = 8'b00110000; assign Signal[2][104] = 8'b00110000; 
assign Signal[0][105] = 8'b01100101; assign Signal[1][105] = 8'b00110001; assign Signal[2][105] = 8'b00110001; 
assign Signal[0][106] = 8'b01100100; assign Signal[1][106] = 8'b00110010; assign Signal[2][106] = 8'b00110010; 
assign Signal[0][107] = 8'b01100011; assign Signal[1][107] = 8'b00110011; assign Signal[2][107] = 8'b00110011; 
assign Signal[0][108] = 8'b01100010; assign Signal[1][108] = 8'b00110100; assign Signal[2][108] = 8'b00110100; 
assign Signal[0][109] = 8'b01100001; assign Signal[1][109] = 8'b00110101; assign Signal[2][109] = 8'b00110101; 
assign Signal[0][110] = 8'b01100000; assign Signal[1][110] = 8'b00110110; assign Signal[2][110] = 8'b00110110; 
assign Signal[0][111] = 8'b01011111; assign Signal[1][111] = 8'b00110111; assign Signal[2][111] = 8'b00110111; 
assign Signal[0][112] = 8'b01011110; assign Signal[1][112] = 8'b00111000; assign Signal[2][112] = 8'b00111000; 
assign Signal[0][113] = 8'b01011100; assign Signal[1][113] = 8'b00111001; assign Signal[2][113] = 8'b00111001; 
assign Signal[0][114] = 8'b01011011; assign Signal[1][114] = 8'b00111010; assign Signal[2][114] = 8'b00111010; 
assign Signal[0][115] = 8'b01011010; assign Signal[1][115] = 8'b00111011; assign Signal[2][115] = 8'b00111011; 
assign Signal[0][116] = 8'b01011001; assign Signal[1][116] = 8'b00111100; assign Signal[2][116] = 8'b00111100; 
assign Signal[0][117] = 8'b01011000; assign Signal[1][117] = 8'b00111101; assign Signal[2][117] = 8'b00111101; 
assign Signal[0][118] = 8'b01010111; assign Signal[1][118] = 8'b00111110; assign Signal[2][118] = 8'b00111110; 
assign Signal[0][119] = 8'b01010101; assign Signal[1][119] = 8'b01000000; assign Signal[2][119] = 8'b01000000; 
assign Signal[0][120] = 8'b01010100; assign Signal[1][120] = 8'b01000001; assign Signal[2][120] = 8'b01000001; 
assign Signal[0][121] = 8'b01010011; assign Signal[1][121] = 8'b01000010; assign Signal[2][121] = 8'b01000010; 
assign Signal[0][122] = 8'b01010010; assign Signal[1][122] = 8'b01000011; assign Signal[2][122] = 8'b01000011; 
assign Signal[0][123] = 8'b01010001; assign Signal[1][123] = 8'b01000100; assign Signal[2][123] = 8'b01000100; 
assign Signal[0][124] = 8'b01001111; assign Signal[1][124] = 8'b01000110; assign Signal[2][124] = 8'b01000110; 
assign Signal[0][125] = 8'b01001110; assign Signal[1][125] = 8'b01000111; assign Signal[2][125] = 8'b01000111; 
assign Signal[0][126] = 8'b01001101; assign Signal[1][126] = 8'b01001000; assign Signal[2][126] = 8'b01001000; 
assign Signal[0][127] = 8'b01001100; assign Signal[1][127] = 8'b01001001; assign Signal[2][127] = 8'b01001001; 
assign Signal[0][128] = 8'b01001011; assign Signal[1][128] = 8'b01001011; assign Signal[2][128] = 8'b01001011; 
assign Signal[0][129] = 8'b01001001; assign Signal[1][129] = 8'b01001100; assign Signal[2][129] = 8'b01001100; 
assign Signal[0][130] = 8'b01001000; assign Signal[1][130] = 8'b01001101; assign Signal[2][130] = 8'b01001101; 
assign Signal[0][131] = 8'b01000111; assign Signal[1][131] = 8'b01001110; assign Signal[2][131] = 8'b01001110; 
assign Signal[0][132] = 8'b01000110; assign Signal[1][132] = 8'b01001111; assign Signal[2][132] = 8'b01001111; 
assign Signal[0][133] = 8'b01000100; assign Signal[1][133] = 8'b01010001; assign Signal[2][133] = 8'b01010001; 
assign Signal[0][134] = 8'b01000011; assign Signal[1][134] = 8'b01010010; assign Signal[2][134] = 8'b01010010; 
assign Signal[0][135] = 8'b01000010; assign Signal[1][135] = 8'b01010011; assign Signal[2][135] = 8'b01010011; 
assign Signal[0][136] = 8'b01000001; assign Signal[1][136] = 8'b01010100; assign Signal[2][136] = 8'b01010100; 
assign Signal[0][137] = 8'b01000000; assign Signal[1][137] = 8'b01010101; assign Signal[2][137] = 8'b01010101; 
assign Signal[0][138] = 8'b00111110; assign Signal[1][138] = 8'b01010111; assign Signal[2][138] = 8'b01010111; 
assign Signal[0][139] = 8'b00111101; assign Signal[1][139] = 8'b01011000; assign Signal[2][139] = 8'b01011000; 
assign Signal[0][140] = 8'b00111100; assign Signal[1][140] = 8'b01011001; assign Signal[2][140] = 8'b01011001; 
assign Signal[0][141] = 8'b00111011; assign Signal[1][141] = 8'b01011010; assign Signal[2][141] = 8'b01011010; 
assign Signal[0][142] = 8'b00111010; assign Signal[1][142] = 8'b01011011; assign Signal[2][142] = 8'b01011011; 
assign Signal[0][143] = 8'b00111001; assign Signal[1][143] = 8'b01011100; assign Signal[2][143] = 8'b01011100; 
assign Signal[0][144] = 8'b00110111; assign Signal[1][144] = 8'b01011101; assign Signal[2][144] = 8'b01011101; 
assign Signal[0][145] = 8'b00110110; assign Signal[1][145] = 8'b01011110; assign Signal[2][145] = 8'b01011110; 
assign Signal[0][146] = 8'b00110101; assign Signal[1][146] = 8'b01011111; assign Signal[2][146] = 8'b01011111; 
assign Signal[0][147] = 8'b00110100; assign Signal[1][147] = 8'b01100000; assign Signal[2][147] = 8'b01100000; 
assign Signal[0][148] = 8'b00110011; assign Signal[1][148] = 8'b01100001; assign Signal[2][148] = 8'b01100001; 
assign Signal[0][149] = 8'b00110010; assign Signal[1][149] = 8'b01100010; assign Signal[2][149] = 8'b01100010; 
assign Signal[0][150] = 8'b00110001; assign Signal[1][150] = 8'b01100011; assign Signal[2][150] = 8'b01100011; 
assign Signal[0][151] = 8'b00110000; assign Signal[1][151] = 8'b01100100; assign Signal[2][151] = 8'b01100100; 
assign Signal[0][152] = 8'b00101111; assign Signal[1][152] = 8'b01100101; assign Signal[2][152] = 8'b01100101; 
assign Signal[0][153] = 8'b00101110; assign Signal[1][153] = 8'b01100110; assign Signal[2][153] = 8'b01100110; 
assign Signal[0][154] = 8'b00101101; assign Signal[1][154] = 8'b01100111; assign Signal[2][154] = 8'b01100111; 
assign Signal[0][155] = 8'b00101100; assign Signal[1][155] = 8'b01101000; assign Signal[2][155] = 8'b01101000; 
assign Signal[0][156] = 8'b00101011; assign Signal[1][156] = 8'b01101001; assign Signal[2][156] = 8'b01101000; 
assign Signal[0][157] = 8'b00101010; assign Signal[1][157] = 8'b01101001; assign Signal[2][157] = 8'b01101001; 
assign Signal[0][158] = 8'b00101001; assign Signal[1][158] = 8'b01101010; assign Signal[2][158] = 8'b01101010; 
assign Signal[0][159] = 8'b00101000; assign Signal[1][159] = 8'b01101011; assign Signal[2][159] = 8'b01101011; 
assign Signal[0][160] = 8'b00100111; assign Signal[1][160] = 8'b01101100; assign Signal[2][160] = 8'b01101011; 
assign Signal[0][161] = 8'b00100110; assign Signal[1][161] = 8'b01101101; assign Signal[2][161] = 8'b01101100; 
assign Signal[0][162] = 8'b00100101; assign Signal[1][162] = 8'b01101101; assign Signal[2][162] = 8'b01101101; 
assign Signal[0][163] = 8'b00100101; assign Signal[1][163] = 8'b01101110; assign Signal[2][163] = 8'b01101101; 
assign Signal[0][164] = 8'b00100100; assign Signal[1][164] = 8'b01101111; assign Signal[2][164] = 8'b01101110; 
assign Signal[0][165] = 8'b00100011; assign Signal[1][165] = 8'b01101111; assign Signal[2][165] = 8'b01101111; 
assign Signal[0][166] = 8'b00100010; assign Signal[1][166] = 8'b01110000; assign Signal[2][166] = 8'b01101111; 
assign Signal[0][167] = 8'b00100010; assign Signal[1][167] = 8'b01110001; assign Signal[2][167] = 8'b01110000; 
assign Signal[0][168] = 8'b00100001; assign Signal[1][168] = 8'b01110001; assign Signal[2][168] = 8'b01110000; 
assign Signal[0][169] = 8'b00100000; assign Signal[1][169] = 8'b01110010; assign Signal[2][169] = 8'b01110001; 
assign Signal[0][170] = 8'b00100000; assign Signal[1][170] = 8'b01110011; assign Signal[2][170] = 8'b01110001; 
assign Signal[0][171] = 8'b00011111; assign Signal[1][171] = 8'b01110011; assign Signal[2][171] = 8'b01110010; 
assign Signal[0][172] = 8'b00011110; assign Signal[1][172] = 8'b01110100; assign Signal[2][172] = 8'b01110010; 
assign Signal[0][173] = 8'b00011110; assign Signal[1][173] = 8'b01110100; assign Signal[2][173] = 8'b01110011; 
assign Signal[0][174] = 8'b00011101; assign Signal[1][174] = 8'b01110101; assign Signal[2][174] = 8'b01110011; 
assign Signal[0][175] = 8'b00011101; assign Signal[1][175] = 8'b01110101; assign Signal[2][175] = 8'b01110011; 
assign Signal[0][176] = 8'b00011100; assign Signal[1][176] = 8'b01110110; assign Signal[2][176] = 8'b01110100; 
assign Signal[0][177] = 8'b00011100; assign Signal[1][177] = 8'b01110110; assign Signal[2][177] = 8'b01110100; 
assign Signal[0][178] = 8'b00011011; assign Signal[1][178] = 8'b01110111; assign Signal[2][178] = 8'b01110101; 
assign Signal[0][179] = 8'b00011011; assign Signal[1][179] = 8'b01110111; assign Signal[2][179] = 8'b01110101; 
assign Signal[0][180] = 8'b00011011; assign Signal[1][180] = 8'b01111000; assign Signal[2][180] = 8'b01110101; 
assign Signal[0][181] = 8'b00011010; assign Signal[1][181] = 8'b01111000; assign Signal[2][181] = 8'b01110110; 
assign Signal[0][182] = 8'b00011010; assign Signal[1][182] = 8'b01111001; assign Signal[2][182] = 8'b01110110; 
assign Signal[0][183] = 8'b00011010; assign Signal[1][183] = 8'b01111001; assign Signal[2][183] = 8'b01110110; 
assign Signal[0][184] = 8'b00011001; assign Signal[1][184] = 8'b01111010; assign Signal[2][184] = 8'b01110110; 
assign Signal[0][185] = 8'b00011001; assign Signal[1][185] = 8'b01111010; assign Signal[2][185] = 8'b01110111; 
assign Signal[0][186] = 8'b00011001; assign Signal[1][186] = 8'b01111010; assign Signal[2][186] = 8'b01110111; 
assign Signal[0][187] = 8'b00011001; assign Signal[1][187] = 8'b01111011; assign Signal[2][187] = 8'b01110111; 
assign Signal[0][188] = 8'b00011001; assign Signal[1][188] = 8'b01111011; assign Signal[2][188] = 8'b01111000; 
assign Signal[0][189] = 8'b00011001; assign Signal[1][189] = 8'b01111100; assign Signal[2][189] = 8'b01111000; 
assign Signal[0][190] = 8'b00011001; assign Signal[1][190] = 8'b01111100; assign Signal[2][190] = 8'b01111000; 
assign Signal[0][191] = 8'b00011001; assign Signal[1][191] = 8'b01111100; assign Signal[2][191] = 8'b01111000; 
assign Signal[0][192] = 8'b00011001; assign Signal[1][192] = 8'b01111101; assign Signal[2][192] = 8'b01111000; 
assign Signal[0][193] = 8'b00011001; assign Signal[1][193] = 8'b01111101; assign Signal[2][193] = 8'b01111001; 
assign Signal[0][194] = 8'b00011001; assign Signal[1][194] = 8'b01111101; assign Signal[2][194] = 8'b01111001; 
assign Signal[0][195] = 8'b00011001; assign Signal[1][195] = 8'b01111110; assign Signal[2][195] = 8'b01111001; 
assign Signal[0][196] = 8'b00011001; assign Signal[1][196] = 8'b01111110; assign Signal[2][196] = 8'b01111001; 
assign Signal[0][197] = 8'b00011001; assign Signal[1][197] = 8'b01111110; assign Signal[2][197] = 8'b01111001; 
assign Signal[0][198] = 8'b00011001; assign Signal[1][198] = 8'b01111111; assign Signal[2][198] = 8'b01111001; 
assign Signal[0][199] = 8'b00011001; assign Signal[1][199] = 8'b01111111; assign Signal[2][199] = 8'b01111010; 
assign Signal[0][200] = 8'b00011001; assign Signal[1][200] = 8'b01111111; assign Signal[2][200] = 8'b01111010; 
assign Signal[0][201] = 8'b00011010; assign Signal[1][201] = 8'b10000000; assign Signal[2][201] = 8'b01111010; 
assign Signal[0][202] = 8'b00011010; assign Signal[1][202] = 8'b10000000; assign Signal[2][202] = 8'b01111010; 
assign Signal[0][203] = 8'b00011010; assign Signal[1][203] = 8'b10000000; assign Signal[2][203] = 8'b01111010; 
assign Signal[0][204] = 8'b00011011; assign Signal[1][204] = 8'b10000000; assign Signal[2][204] = 8'b01111010; 
assign Signal[0][205] = 8'b00011011; assign Signal[1][205] = 8'b10000001; assign Signal[2][205] = 8'b01111010; 
assign Signal[0][206] = 8'b00011011; assign Signal[1][206] = 8'b10000001; assign Signal[2][206] = 8'b01111010; 
assign Signal[0][207] = 8'b00011100; assign Signal[1][207] = 8'b10000001; assign Signal[2][207] = 8'b01111010; 
assign Signal[0][208] = 8'b00011100; assign Signal[1][208] = 8'b10000001; assign Signal[2][208] = 8'b01111011; 
assign Signal[0][209] = 8'b00011101; assign Signal[1][209] = 8'b10000010; assign Signal[2][209] = 8'b01111011; 
assign Signal[0][210] = 8'b00011101; assign Signal[1][210] = 8'b10000010; assign Signal[2][210] = 8'b01111011; 
assign Signal[0][211] = 8'b00011110; assign Signal[1][211] = 8'b10000010; assign Signal[2][211] = 8'b01111011; 
assign Signal[0][212] = 8'b00011110; assign Signal[1][212] = 8'b10000010; assign Signal[2][212] = 8'b01111011; 
assign Signal[0][213] = 8'b00011111; assign Signal[1][213] = 8'b10000011; assign Signal[2][213] = 8'b01111011; 
assign Signal[0][214] = 8'b00100000; assign Signal[1][214] = 8'b10000011; assign Signal[2][214] = 8'b01111011; 
assign Signal[0][215] = 8'b00100000; assign Signal[1][215] = 8'b10000011; assign Signal[2][215] = 8'b01111011; 
assign Signal[0][216] = 8'b00100001; assign Signal[1][216] = 8'b10000011; assign Signal[2][216] = 8'b01111011; 
assign Signal[0][217] = 8'b00100010; assign Signal[1][217] = 8'b10000100; assign Signal[2][217] = 8'b01111011; 
assign Signal[0][218] = 8'b00100010; assign Signal[1][218] = 8'b10000100; assign Signal[2][218] = 8'b01111011; 
assign Signal[0][219] = 8'b00100011; assign Signal[1][219] = 8'b10000100; assign Signal[2][219] = 8'b01111011; 
assign Signal[0][220] = 8'b00100100; assign Signal[1][220] = 8'b10000100; assign Signal[2][220] = 8'b01111011; 
assign Signal[0][221] = 8'b00100101; assign Signal[1][221] = 8'b10000100; assign Signal[2][221] = 8'b01111011; 
assign Signal[0][222] = 8'b00100101; assign Signal[1][222] = 8'b10000101; assign Signal[2][222] = 8'b01111100; 
assign Signal[0][223] = 8'b00100110; assign Signal[1][223] = 8'b10000101; assign Signal[2][223] = 8'b01111100; 
assign Signal[0][224] = 8'b00100111; assign Signal[1][224] = 8'b10000101; assign Signal[2][224] = 8'b01111100; 
assign Signal[0][225] = 8'b00101000; assign Signal[1][225] = 8'b10000101; assign Signal[2][225] = 8'b01111100; 
assign Signal[0][226] = 8'b00101001; assign Signal[1][226] = 8'b10000101; assign Signal[2][226] = 8'b01111100; 
assign Signal[0][227] = 8'b00101010; assign Signal[1][227] = 8'b10000110; assign Signal[2][227] = 8'b01111100; 
assign Signal[0][228] = 8'b00101011; assign Signal[1][228] = 8'b10000110; assign Signal[2][228] = 8'b01111100; 
assign Signal[0][229] = 8'b00101100; assign Signal[1][229] = 8'b10000110; assign Signal[2][229] = 8'b01111100; 
assign Signal[0][230] = 8'b00101101; assign Signal[1][230] = 8'b10000110; assign Signal[2][230] = 8'b01111100; 
assign Signal[0][231] = 8'b00101110; assign Signal[1][231] = 8'b10000110; assign Signal[2][231] = 8'b01111100; 
assign Signal[0][232] = 8'b00101111; assign Signal[1][232] = 8'b10000110; assign Signal[2][232] = 8'b01111100; 
assign Signal[0][233] = 8'b00110000; assign Signal[1][233] = 8'b10000111; assign Signal[2][233] = 8'b01111100; 
assign Signal[0][234] = 8'b00110001; assign Signal[1][234] = 8'b10000111; assign Signal[2][234] = 8'b01111100; 
assign Signal[0][235] = 8'b00110010; assign Signal[1][235] = 8'b10000111; assign Signal[2][235] = 8'b01111100; 
assign Signal[0][236] = 8'b00110011; assign Signal[1][236] = 8'b10000111; assign Signal[2][236] = 8'b01111100; 
assign Signal[0][237] = 8'b00110100; assign Signal[1][237] = 8'b10000111; assign Signal[2][237] = 8'b01111100; 
assign Signal[0][238] = 8'b00110101; assign Signal[1][238] = 8'b10000111; assign Signal[2][238] = 8'b01111100; 
assign Signal[0][239] = 8'b00110110; assign Signal[1][239] = 8'b10000111; assign Signal[2][239] = 8'b01111100; 
assign Signal[0][240] = 8'b00110111; assign Signal[1][240] = 8'b10001000; assign Signal[2][240] = 8'b01111100; 
assign Signal[0][241] = 8'b00111001; assign Signal[1][241] = 8'b10001000; assign Signal[2][241] = 8'b01111100; 
assign Signal[0][242] = 8'b00111010; assign Signal[1][242] = 8'b10001000; assign Signal[2][242] = 8'b01111100; 
assign Signal[0][243] = 8'b00111011; assign Signal[1][243] = 8'b10001000; assign Signal[2][243] = 8'b01111100; 
assign Signal[0][244] = 8'b00111100; assign Signal[1][244] = 8'b10001000; assign Signal[2][244] = 8'b01111100; 
assign Signal[0][245] = 8'b00111101; assign Signal[1][245] = 8'b10001000; assign Signal[2][245] = 8'b01111100; 
assign Signal[0][246] = 8'b00111110; assign Signal[1][246] = 8'b10001000; assign Signal[2][246] = 8'b01111100; 
assign Signal[0][247] = 8'b01000000; assign Signal[1][247] = 8'b10001001; assign Signal[2][247] = 8'b01111100; 
assign Signal[0][248] = 8'b01000001; assign Signal[1][248] = 8'b10001001; assign Signal[2][248] = 8'b01111100; 
assign Signal[0][249] = 8'b01000010; assign Signal[1][249] = 8'b10001001; assign Signal[2][249] = 8'b01111100; 
assign Signal[0][250] = 8'b01000011; assign Signal[1][250] = 8'b10001001; assign Signal[2][250] = 8'b01111100; 
assign Signal[0][251] = 8'b01000100; assign Signal[1][251] = 8'b10001001; assign Signal[2][251] = 8'b01111100; 
assign Signal[0][252] = 8'b01000110; assign Signal[1][252] = 8'b10001001; assign Signal[2][252] = 8'b01111100; 
assign Signal[0][253] = 8'b01000111; assign Signal[1][253] = 8'b10001001; assign Signal[2][253] = 8'b01111100; 
assign Signal[0][254] = 8'b01001000; assign Signal[1][254] = 8'b10001001; assign Signal[2][254] = 8'b01111100; 
assign Signal[0][255] = 8'b01001001; assign Signal[1][255] = 8'b10001010; assign Signal[2][255] = 8'b01111100; 


*/

  /* Sequential Logic */
  always @(negedge clk) begin
    busy_counter <= busy_counter +1'b1;
    if (busy_counter == SIZE_b) begin
    addr <= addr + 1'b1;
    signal_q <= Signal [0][addr];
    //signal_q <= addr;
    end 
  end
  
// Try an innitial block here for just loading in all the values to read only memory.   


initial begin // sets all initial values to 0. 
 Signal[0][0] <= 8'b01001011;  Signal[1][0] <= 8'b00001011;  Signal[2][0] <= 8'b00000000; 
 Signal[0][1] <= 8'b01001100;  Signal[1][1] <= 8'b00001011;  Signal[2][1] <= 8'b00000000; 
 Signal[0][2] <= 8'b01001101;  Signal[1][2] <= 8'b00001100;  Signal[2][2] <= 8'b00000000; 
 Signal[0][3] <= 8'b01001110;  Signal[1][3] <= 8'b00001100;  Signal[2][3] <= 8'b00000000; 
 Signal[0][4] <= 8'b01001111;  Signal[1][4] <= 8'b00001100;  Signal[2][4] <= 8'b00000000; 
 Signal[0][5] <= 8'b01010001;  Signal[1][5] <= 8'b00001100;  Signal[2][5] <= 8'b00000000; 
 Signal[0][6] <= 8'b01010010;  Signal[1][6] <= 8'b00001100;  Signal[2][6] <= 8'b00000000; 
 Signal[0][7] <= 8'b01010011;  Signal[1][7] <= 8'b00001100;  Signal[2][7] <= 8'b00000000; 
 Signal[0][8] <= 8'b01010100;  Signal[1][8] <= 8'b00001100;  Signal[2][8] <= 8'b00000000; 
 Signal[0][9] <= 8'b01010101;  Signal[1][9] <= 8'b00001100;  Signal[2][9] <= 8'b00000000; 
 Signal[0][10] <= 8'b01010111;  Signal[1][10] <= 8'b00001101;  Signal[2][10] <= 8'b0; 
 Signal[0][11] <= 8'b01011000;  Signal[1][11] <= 8'b00001101;  Signal[2][11] <= 8'b0; 
 Signal[0][12] <= 8'b01011001;  Signal[1][12] <= 8'b00001101;  Signal[2][12] <= 8'h00; 
 Signal[0][13] <= 8'b01011010;  Signal[1][13] <= 8'b00001101;  Signal[2][13] <= 8'hFF; 
 Signal[0][14] <= 8'b01011011;  Signal[1][14] <= 8'b00001101;  Signal[2][14] <= 8'hFF; 
 Signal[0][15] <= 8'b01011100;  Signal[1][15] <= 8'b00001101;  Signal[2][15] <= 8'b0; 
 Signal[0][16] <= 8'b01011110;  Signal[1][16] <= 8'b00001101;  Signal[2][16] <= 8'b0; 
 Signal[0][17] <= 8'b01011111;  Signal[1][17] <= 8'b00001110;  Signal[2][17] <= 8'b0; 
 Signal[0][18] <= 8'b01100000;  Signal[1][18] <= 8'b00001110;  Signal[2][18] <= 8'b0; 
 Signal[0][19] <= 8'b01100001;  Signal[1][19] <= 8'b00001110;  Signal[2][19] <= 8'b0; 
 Signal[0][20] <= 8'b01100010;  Signal[1][20] <= 8'b00001110;  Signal[2][20] <= 8'b0; 
 Signal[0][21] <= 8'b01100011;  Signal[1][21] <= 8'b00001110;  Signal[2][21] <= 8'b0; 
 Signal[0][22] <= 8'b01100100;  Signal[1][22] <= 8'b00001110;  Signal[2][22] <= 8'b0; 
 Signal[0][23] <= 8'b01100101;  Signal[1][23] <= 8'b00001110;  Signal[2][23] <= 8'b00000000; 
 Signal[0][24] <= 8'b01100110;  Signal[1][24] <= 8'b00001111;  Signal[2][24] <= 8'b00000000; 
 Signal[0][25] <= 8'b01100111;  Signal[1][25] <= 8'b00001111;  Signal[2][25] <= 8'b00000000; 
 Signal[0][26] <= 8'b01101000;  Signal[1][26] <= 8'b00001111;  Signal[2][26] <= 8'b00000000; 
 Signal[0][27] <= 8'b01101001;  Signal[1][27] <= 8'b00001111;  Signal[2][27] <= 8'b00000000; 
 Signal[0][28] <= 8'b01101010;  Signal[1][28] <= 8'b00001111;  Signal[2][28] <= 8'b00000000; 
 Signal[0][29] <= 8'b01101011;  Signal[1][29] <= 8'b00001111;  Signal[2][29] <= 8'b00000000; 
 Signal[0][30] <= 8'b01101100;  Signal[1][30] <= 8'b00010000;  Signal[2][30] <= 8'b00000000; 
 Signal[0][31] <= 8'b01101101;  Signal[1][31] <= 8'b00010000;  Signal[2][31] <= 8'b00000000; 
 Signal[0][32] <= 8'b01101110;  Signal[1][32] <= 8'b00010000;  Signal[2][32] <= 8'b00000000; 
 Signal[0][33] <= 8'b01101111;  Signal[1][33] <= 8'b00010000;  Signal[2][33] <= 8'b00000000; 
 Signal[0][34] <= 8'b01110000;  Signal[1][34] <= 8'b00010000;  Signal[2][34] <= 8'b00000000; 
 Signal[0][35] <= 8'b01110000;  Signal[1][35] <= 8'b00010001;  Signal[2][35] <= 8'b00000000; 
 Signal[0][36] <= 8'b01110001;  Signal[1][36] <= 8'b00010001;  Signal[2][36] <= 8'b00000000; 
 Signal[0][37] <= 8'b01110010;  Signal[1][37] <= 8'b00010001;  Signal[2][37] <= 8'b00000000; 
 Signal[0][38] <= 8'b01110011;  Signal[1][38] <= 8'b00010001;  Signal[2][38] <= 8'b00000000; 
 Signal[0][39] <= 8'b01110011;  Signal[1][39] <= 8'b00010001;  Signal[2][39] <= 8'b00000000; 
 Signal[0][40] <= 8'b01110100;  Signal[1][40] <= 8'b00010010;  Signal[2][40] <= 8'b00000000; 
 Signal[0][41] <= 8'b01110101;  Signal[1][41] <= 8'b00010010;  Signal[2][41] <= 8'b00000000; 
 Signal[0][42] <= 8'b01110101;  Signal[1][42] <= 8'b00010010;  Signal[2][42] <= 8'b00000000; 
 Signal[0][43] <= 8'b01110110;  Signal[1][43] <= 8'b00010010;  Signal[2][43] <= 8'b00000000; 
 Signal[0][44] <= 8'b01110111;  Signal[1][44] <= 8'b00010011;  Signal[2][44] <= 8'b00000000; 
 Signal[0][45] <= 8'b01110111;  Signal[1][45] <= 8'b00010011;  Signal[2][45] <= 8'b00000000; 
 Signal[0][46] <= 8'b01111000;  Signal[1][46] <= 8'b00010011;  Signal[2][46] <= 8'b00000000; 
 Signal[0][47] <= 8'b01111000;  Signal[1][47] <= 8'b00010011;  Signal[2][47] <= 8'b00000000; 
 Signal[0][48] <= 8'b01111001;  Signal[1][48] <= 8'b00010100;  Signal[2][48] <= 8'b00000000; 
 Signal[0][49] <= 8'b01111001;  Signal[1][49] <= 8'b00010100;  Signal[2][49] <= 8'b00000000; 
 Signal[0][50] <= 8'b01111010;  Signal[1][50] <= 8'b00010100;  Signal[2][50] <= 8'b00000000; 
 Signal[0][51] <= 8'b01111010;  Signal[1][51] <= 8'b00010100;  Signal[2][51] <= 8'b00000000; 
 Signal[0][52] <= 8'b01111010;  Signal[1][52] <= 8'b00010101;  Signal[2][52] <= 8'b00000000; 
 Signal[0][53] <= 8'b01111011;  Signal[1][53] <= 8'b00010101;  Signal[2][53] <= 8'b00000000; 
 Signal[0][54] <= 8'b01111011;  Signal[1][54] <= 8'b00010101;  Signal[2][54] <= 8'b00000000; 
 Signal[0][55] <= 8'b01111011;  Signal[1][55] <= 8'b00010101;  Signal[2][55] <= 8'b00000000; 
 Signal[0][56] <= 8'b01111100;  Signal[1][56] <= 8'b00010110;  Signal[2][56] <= 8'b00000000; 
 Signal[0][57] <= 8'b01111100;  Signal[1][57] <= 8'b00010110;  Signal[2][57] <= 8'b00000000; 
 Signal[0][58] <= 8'b01111100;  Signal[1][58] <= 8'b00010110;  Signal[2][58] <= 8'b00000000; 
 Signal[0][59] <= 8'b01111100;  Signal[1][59] <= 8'b00010111;  Signal[2][59] <= 8'b00000000; 
 Signal[0][60] <= 8'b01111100;  Signal[1][60] <= 8'b00010111;  Signal[2][60] <= 8'b00000000; 
 Signal[0][61] <= 8'b01111100;  Signal[1][61] <= 8'b00010111;  Signal[2][61] <= 8'b00000000; 
 Signal[0][62] <= 8'b01111100;  Signal[1][62] <= 8'b00011000;  Signal[2][62] <= 8'b00000000; 
 Signal[0][63] <= 8'b01111100;  Signal[1][63] <= 8'b00011000;  Signal[2][63] <= 8'b00000000; 
 Signal[0][64] <= 8'b01111101;  Signal[1][64] <= 8'b00011000;  Signal[2][64] <= 8'b00000000; 
 Signal[0][65] <= 8'b01111100;  Signal[1][65] <= 8'b00011001;  Signal[2][65] <= 8'b00000000; 
 Signal[0][66] <= 8'b01111100;  Signal[1][66] <= 8'b00011001;  Signal[2][66] <= 8'b00000000; 
 Signal[0][67] <= 8'b01111100;  Signal[1][67] <= 8'b00011001;  Signal[2][67] <= 8'b00000000; 
 Signal[0][68] <= 8'b01111100;  Signal[1][68] <= 8'b00011010;  Signal[2][68] <= 8'b00000000; 
 Signal[0][69] <= 8'b01111100;  Signal[1][69] <= 8'b00011010;  Signal[2][69] <= 8'b00000000; 
 Signal[0][70] <= 8'b01111100;  Signal[1][70] <= 8'b00011011;  Signal[2][70] <= 8'b00000000; 
 Signal[0][71] <= 8'b01111100;  Signal[1][71] <= 8'b00011011;  Signal[2][71] <= 8'b00000000; 
 Signal[0][72] <= 8'b01111100;  Signal[1][72] <= 8'b00011011;  Signal[2][72] <= 8'b00000000; 
 Signal[0][73] <= 8'b01111011;  Signal[1][73] <= 8'b00011100;  Signal[2][73] <= 8'b00000000; 
 Signal[0][74] <= 8'b01111011;  Signal[1][74] <= 8'b00011100;  Signal[2][74] <= 8'b00000000; 
 Signal[0][75] <= 8'b01111011;  Signal[1][75] <= 8'b00011101;  Signal[2][75] <= 8'b00000000; 
 Signal[0][76] <= 8'b01111010;  Signal[1][76] <= 8'b00011101;  Signal[2][76] <= 8'b00000000; 
 Signal[0][77] <= 8'b01111010;  Signal[1][77] <= 8'b00011110;  Signal[2][77] <= 8'b00000000; 
 Signal[0][78] <= 8'b01111010;  Signal[1][78] <= 8'b00011110;  Signal[2][78] <= 8'b00000000; 
 Signal[0][79] <= 8'b01111001;  Signal[1][79] <= 8'b00011111;  Signal[2][79] <= 8'b00000000; 
 Signal[0][80] <= 8'b01111001;  Signal[1][80] <= 8'b00011111;  Signal[2][80] <= 8'b00000000; 
 Signal[0][81] <= 8'b01111000;  Signal[1][81] <= 8'b00100000;  Signal[2][81] <= 8'b00000000; 
 Signal[0][82] <= 8'b01111000;  Signal[1][82] <= 8'b00100000;  Signal[2][82] <= 8'b00000000; 
 Signal[0][83] <= 8'b01110111;  Signal[1][83] <= 8'b00100001;  Signal[2][83] <= 8'b00000000; 
 Signal[0][84] <= 8'b01110111;  Signal[1][84] <= 8'b00100001;  Signal[2][84] <= 8'b00000000; 
 Signal[0][85] <= 8'b01110110;  Signal[1][85] <= 8'b00100010;  Signal[2][85] <= 8'b00000000; 
 Signal[0][86] <= 8'b01110101;  Signal[1][86] <= 8'b00100010;  Signal[2][86] <= 8'b00000000; 
 Signal[0][87] <= 8'b01110101;  Signal[1][87] <= 8'b00100011;  Signal[2][87] <= 8'b00000000; 
 Signal[0][88] <= 8'b01110100;  Signal[1][88] <= 8'b00100100;  Signal[2][88] <= 8'b00000000; 
 Signal[0][89] <= 8'b01110011;  Signal[1][89] <= 8'b00100100;  Signal[2][89] <= 8'b00000000; 
 Signal[0][90] <= 8'b01110011;  Signal[1][90] <= 8'b00100101;  Signal[2][90] <= 8'b00000000; 
 Signal[0][91] <= 8'b01110010;  Signal[1][91] <= 8'b00100110;  Signal[2][91] <= 8'b00000000; 
 Signal[0][92] <= 8'b01110001;  Signal[1][92] <= 8'b00100110;  Signal[2][92] <= 8'b00000000; 
 Signal[0][93] <= 8'b01110000;  Signal[1][93] <= 8'b00100111;  Signal[2][93] <= 8'b00000000; 
 Signal[0][94] <= 8'b01110000;  Signal[1][94] <= 8'b00101000;  Signal[2][94] <= 8'b00000000; 
 Signal[0][95] <= 8'b01101111;  Signal[1][95] <= 8'b00101000;  Signal[2][95] <= 8'b00000000; 
 Signal[0][96] <= 8'b01101110;  Signal[1][96] <= 8'b00101001;  Signal[2][96] <= 8'b00000000; 
 Signal[0][97] <= 8'b01101101;  Signal[1][97] <= 8'b00101010;  Signal[2][97] <= 8'b00000000; 
 Signal[0][98] <= 8'b01101100;  Signal[1][98] <= 8'b00101011;  Signal[2][98] <= 8'b00000000; 
 Signal[0][99] <= 8'b01101011;  Signal[1][99] <= 8'b00101100;  Signal[2][99] <= 8'b00000000; 
 Signal[0][100] <= 8'b01101010;  Signal[1][100] <= 8'b00101100;  Signal[2][100] <= 8'b00000000; 
 Signal[0][101] <= 8'b01101001;  Signal[1][101] <= 8'b00101101;  Signal[2][101] <= 8'b00000000; 
 Signal[0][102] <= 8'b01101000;  Signal[1][102] <= 8'b00101110;  Signal[2][102] <= 8'b00000000; 
 Signal[0][103] <= 8'b01100111;  Signal[1][103] <= 8'b00101111;  Signal[2][103] <= 8'b00000000; 
 Signal[0][104] <= 8'b01100110;  Signal[1][104] <= 8'b00110000;  Signal[2][104] <= 8'b00000000; 
 Signal[0][105] <= 8'b01100101;  Signal[1][105] <= 8'b00110001;  Signal[2][105] <= 8'b00000000; 
 Signal[0][106] <= 8'b01100100;  Signal[1][106] <= 8'b00110010;  Signal[2][106] <= 8'b00000000; 
 Signal[0][107] <= 8'b01100011;  Signal[1][107] <= 8'b00110011;  Signal[2][107] <= 8'b00000000; 
 Signal[0][108] <= 8'b01100010;  Signal[1][108] <= 8'b00110100;  Signal[2][108] <= 8'b00000000; 
 Signal[0][109] <= 8'b01100001;  Signal[1][109] <= 8'b00110101;  Signal[2][109] <= 8'b00000000; 
 Signal[0][110] <= 8'b01100000;  Signal[1][110] <= 8'b00110110;  Signal[2][110] <= 8'b00000000; 
 Signal[0][111] <= 8'b01011111;  Signal[1][111] <= 8'b00110111;  Signal[2][111] <= 8'b00000000; 
 Signal[0][112] <= 8'b01011110;  Signal[1][112] <= 8'b00111000;  Signal[2][112] <= 8'b00000000; 
 Signal[0][113] <= 8'b01011100;  Signal[1][113] <= 8'b00111001;  Signal[2][113] <= 8'b00000000; 
 Signal[0][114] <= 8'b01011011;  Signal[1][114] <= 8'b00111010;  Signal[2][114] <= 8'b00000000; 
 Signal[0][115] <= 8'b01011010;  Signal[1][115] <= 8'b00111011;  Signal[2][115] <= 8'b00000000; 
 Signal[0][116] <= 8'b01011001;  Signal[1][116] <= 8'b00111100;  Signal[2][116] <= 8'b00000000; 
 Signal[0][117] <= 8'b01011000;  Signal[1][117] <= 8'b00111101;  Signal[2][117] <= 8'b00000000; 
 Signal[0][118] <= 8'b01010111;  Signal[1][118] <= 8'b00111110;  Signal[2][118] <= 8'b00000000; 
 Signal[0][119] <= 8'b01010101;  Signal[1][119] <= 8'b01000000;  Signal[2][119] <= 8'b00000000; 
 Signal[0][120] <= 8'b01010100;  Signal[1][120] <= 8'b01000001;  Signal[2][120] <= 8'b00000000; 
 Signal[0][121] <= 8'b01010011;  Signal[1][121] <= 8'b01000010;  Signal[2][121] <= 8'b00000000; 
 Signal[0][122] <= 8'b01010010;  Signal[1][122] <= 8'b01000011;  Signal[2][122] <= 8'b00000000; 
 Signal[0][123] <= 8'b01010001;  Signal[1][123] <= 8'b01000100;  Signal[2][123] <= 8'b00000000; 
 Signal[0][124] <= 8'b01001111;  Signal[1][124] <= 8'b01000110;  Signal[2][124] <= 8'b00000000; 
 Signal[0][125] <= 8'b01001110;  Signal[1][125] <= 8'b01000111;  Signal[2][125] <= 8'b00000000; 
 Signal[0][126] <= 8'b01001101;  Signal[1][126] <= 8'b01001000;  Signal[2][126] <= 8'b00000000; 
 Signal[0][127] <= 8'b01001100;  Signal[1][127] <= 8'b01001001;  Signal[2][127] <= 8'b00000000; 
 Signal[0][128] <= 8'b01001011;  Signal[1][128] <= 8'b01001011;  Signal[2][128] <= 8'b00000000; 
 Signal[0][129] <= 8'b01001001;  Signal[1][129] <= 8'b01001100;  Signal[2][129] <= 8'b00000000; 
 Signal[0][130] <= 8'b01001000;  Signal[1][130] <= 8'b01001101;  Signal[2][130] <= 8'b00000000; 
 Signal[0][131] <= 8'b01000111;  Signal[1][131] <= 8'b01001110;  Signal[2][131] <= 8'b00000000; 
 Signal[0][132] <= 8'b01000110;  Signal[1][132] <= 8'b01001111;  Signal[2][132] <= 8'b00000000; 
 Signal[0][133] <= 8'b01000100;  Signal[1][133] <= 8'b01010001;  Signal[2][133] <= 8'b00000000; 
 Signal[0][134] <= 8'b01000011;  Signal[1][134] <= 8'b01010010;  Signal[2][134] <= 8'b00000000; 
 Signal[0][135] <= 8'b01000010;  Signal[1][135] <= 8'b01010011;  Signal[2][135] <= 8'b00000000; 
 Signal[0][136] <= 8'b01000001;  Signal[1][136] <= 8'b01010100;  Signal[2][136] <= 8'b00000000; 
 Signal[0][137] <= 8'b01000000;  Signal[1][137] <= 8'b01010101;  Signal[2][137] <= 8'b00000000; 
 Signal[0][138] <= 8'b00111110;  Signal[1][138] <= 8'b01010111;  Signal[2][138] <= 8'b00000000; 
 Signal[0][139] <= 8'b00111101;  Signal[1][139] <= 8'b01011000;  Signal[2][139] <= 8'b00000000; 
 Signal[0][140] <= 8'b00111100;  Signal[1][140] <= 8'b01011001;  Signal[2][140] <= 8'b00000000; 
 Signal[0][141] <= 8'b00111011;  Signal[1][141] <= 8'b01011010;  Signal[2][141] <= 8'b00000000; 
 Signal[0][142] <= 8'b00111010;  Signal[1][142] <= 8'b01011011;  Signal[2][142] <= 8'b00000000; 
 Signal[0][143] <= 8'b00111001;  Signal[1][143] <= 8'b01011100;  Signal[2][143] <= 8'b00000000; 
 Signal[0][144] <= 8'b00110111;  Signal[1][144] <= 8'b01011101;  Signal[2][144] <= 8'b00000000; 
 Signal[0][145] <= 8'b00110110;  Signal[1][145] <= 8'b01011110;  Signal[2][145] <= 8'b00000000; 
 Signal[0][146] <= 8'b00110101;  Signal[1][146] <= 8'b01011111;  Signal[2][146] <= 8'b00000000; 
 Signal[0][147] <= 8'b00110100;  Signal[1][147] <= 8'b01100000;  Signal[2][147] <= 8'b00000000; 
 Signal[0][148] <= 8'b00110011;  Signal[1][148] <= 8'b01100001;  Signal[2][148] <= 8'b00000000; 
 Signal[0][149] <= 8'b00110010;  Signal[1][149] <= 8'b01100010;  Signal[2][149] <= 8'b00000000; 
 Signal[0][150] <= 8'b00110001;  Signal[1][150] <= 8'b01100011;  Signal[2][150] <= 8'b00000000; 
 Signal[0][151] <= 8'b00110000;  Signal[1][151] <= 8'b01100100;  Signal[2][151] <= 8'b00000000; 
 Signal[0][152] <= 8'b00101111;  Signal[1][152] <= 8'b01100101;  Signal[2][152] <= 8'b00000000; 
 Signal[0][153] <= 8'b00101110;  Signal[1][153] <= 8'b01100110;  Signal[2][153] <= 8'b00000000; 
 Signal[0][154] <= 8'b00101101;  Signal[1][154] <= 8'b01100111;  Signal[2][154] <= 8'b00000000; 
 Signal[0][155] <= 8'b00101100;  Signal[1][155] <= 8'b01101000;  Signal[2][155] <= 8'b00000000; 
 Signal[0][156] <= 8'b00101011;  Signal[1][156] <= 8'b01101001;  Signal[2][156] <= 8'b00000000; 
 Signal[0][157] <= 8'b00101010;  Signal[1][157] <= 8'b01101001;  Signal[2][157] <= 8'b00000000; 
 Signal[0][158] <= 8'b00101001;  Signal[1][158] <= 8'b01101010;  Signal[2][158] <= 8'b00000000; 
 Signal[0][159] <= 8'b00101000;  Signal[1][159] <= 8'b01101011;  Signal[2][159] <= 8'b00000000; 
 Signal[0][160] <= 8'b00100111;  Signal[1][160] <= 8'b01101100;  Signal[2][160] <= 8'b00000000; 
 Signal[0][161] <= 8'b00100110;  Signal[1][161] <= 8'b01101101;  Signal[2][161] <= 8'b00000000; 
 Signal[0][162] <= 8'b00100101;  Signal[1][162] <= 8'b01101101;  Signal[2][162] <= 8'b00000000; 
 Signal[0][163] <= 8'b00100101;  Signal[1][163] <= 8'b01101110;  Signal[2][163] <= 8'b00000000; 
 Signal[0][164] <= 8'b00100100;  Signal[1][164] <= 8'b01101111;  Signal[2][164] <= 8'b00000000; 
 Signal[0][165] <= 8'b00100011;  Signal[1][165] <= 8'b01101111;  Signal[2][165] <= 8'b00000000; 
 Signal[0][166] <= 8'b00100010;  Signal[1][166] <= 8'b01110000;  Signal[2][166] <= 8'b00000000; 
 Signal[0][167] <= 8'b00100010;  Signal[1][167] <= 8'b01110001;  Signal[2][167] <= 8'b00000000; 
 Signal[0][168] <= 8'b00100001;  Signal[1][168] <= 8'b01110001;  Signal[2][168] <= 8'b00000000; 
 Signal[0][169] <= 8'b00100000;  Signal[1][169] <= 8'b01110010;  Signal[2][169] <= 8'b00000000; 
 Signal[0][170] <= 8'b00100000;  Signal[1][170] <= 8'b01110011;  Signal[2][170] <= 8'b00000000; 
 Signal[0][171] <= 8'b00011111;  Signal[1][171] <= 8'b01110011;  Signal[2][171] <= 8'b00000000; 
 Signal[0][172] <= 8'b00011110;  Signal[1][172] <= 8'b01110100;  Signal[2][172] <= 8'b00000000; 
 Signal[0][173] <= 8'b00011110;  Signal[1][173] <= 8'b01110100;  Signal[2][173] <= 8'b00000000; 
 Signal[0][174] <= 8'b00011101;  Signal[1][174] <= 8'b01110101;  Signal[2][174] <= 8'b00000000; 
 Signal[0][175] <= 8'b00011101;  Signal[1][175] <= 8'b01110101;  Signal[2][175] <= 8'b00000000; 
 Signal[0][176] <= 8'b00011100;  Signal[1][176] <= 8'b01110110;  Signal[2][176] <= 8'b00000000; 
 Signal[0][177] <= 8'b00011100;  Signal[1][177] <= 8'b01110110;  Signal[2][177] <= 8'b00000000; 
 Signal[0][178] <= 8'b00011011;  Signal[1][178] <= 8'b01110111;  Signal[2][178] <= 8'b00000000; 
 Signal[0][179] <= 8'b00011011;  Signal[1][179] <= 8'b01110111;  Signal[2][179] <= 8'b00000000; 
 Signal[0][180] <= 8'b00011011;  Signal[1][180] <= 8'b01111000;  Signal[2][180] <= 8'b00000000; 
 Signal[0][181] <= 8'b00011010;  Signal[1][181] <= 8'b01111000;  Signal[2][181] <= 8'b00000000; 
 Signal[0][182] <= 8'b00011010;  Signal[1][182] <= 8'b01111001;  Signal[2][182] <= 8'b00000000; 
 Signal[0][183] <= 8'b00011010;  Signal[1][183] <= 8'b01111001;  Signal[2][183] <= 8'b00000000; 
 Signal[0][184] <= 8'b00011001;  Signal[1][184] <= 8'b01111010;  Signal[2][184] <= 8'b00000000; 
 Signal[0][185] <= 8'b00011001;  Signal[1][185] <= 8'b01111010;  Signal[2][185] <= 8'b00000000; 
 Signal[0][186] <= 8'b00011001;  Signal[1][186] <= 8'b01111010;  Signal[2][186] <= 8'b00000000; 
 Signal[0][187] <= 8'b00011001;  Signal[1][187] <= 8'b01111011;  Signal[2][187] <= 8'b00000000; 
 Signal[0][188] <= 8'b00011001;  Signal[1][188] <= 8'b01111011;  Signal[2][188] <= 8'b00000000; 
 Signal[0][189] <= 8'b00011001;  Signal[1][189] <= 8'b01111100;  Signal[2][189] <= 8'b00000000; 
 Signal[0][190] <= 8'b00011001;  Signal[1][190] <= 8'b01111100;  Signal[2][190] <= 8'b00000000; 
 Signal[0][191] <= 8'b00011001;  Signal[1][191] <= 8'b01111100;  Signal[2][191] <= 8'b00000000; 
 Signal[0][192] <= 8'b00011001;  Signal[1][192] <= 8'b01111101;  Signal[2][192] <= 8'b00000000; 
 Signal[0][193] <= 8'b00011001;  Signal[1][193] <= 8'b01111101;  Signal[2][193] <= 8'b00000000; 
 Signal[0][194] <= 8'b00011001;  Signal[1][194] <= 8'b01111101;  Signal[2][194] <= 8'b00000000; 
 Signal[0][195] <= 8'b00011001;  Signal[1][195] <= 8'b01111110;  Signal[2][195] <= 8'b00000000; 
 Signal[0][196] <= 8'b00011001;  Signal[1][196] <= 8'b01111110;  Signal[2][196] <= 8'b00000000; 
 Signal[0][197] <= 8'b00011001;  Signal[1][197] <= 8'b01111110;  Signal[2][197] <= 8'b00000000; 
 Signal[0][198] <= 8'b00011001;  Signal[1][198] <= 8'b01111111;  Signal[2][198] <= 8'b00000000; 
 Signal[0][199] <= 8'b00011001;  Signal[1][199] <= 8'b01111111;  Signal[2][199] <= 8'b00000000; 
 Signal[0][200] <= 8'b00011001;  Signal[1][200] <= 8'b01111111;  Signal[2][200] <= 8'b00000000; 
 Signal[0][201] <= 8'b00011010;  Signal[1][201] <= 8'b10000000;  Signal[2][201] <= 8'b00000000; 
 Signal[0][202] <= 8'b00011010;  Signal[1][202] <= 8'b10000000;  Signal[2][202] <= 8'b00000000; 
 Signal[0][203] <= 8'b00011010;  Signal[1][203] <= 8'b10000000;  Signal[2][203] <= 8'b00000000; 
 Signal[0][204] <= 8'b00011011;  Signal[1][204] <= 8'b10000000;  Signal[2][204] <= 8'b00000000; 
 Signal[0][205] <= 8'b00011011;  Signal[1][205] <= 8'b10000001;  Signal[2][205] <= 8'b00000000; 
 Signal[0][206] <= 8'b00011011;  Signal[1][206] <= 8'b10000001;  Signal[2][206] <= 8'b00000000; 
 Signal[0][207] <= 8'b00011100;  Signal[1][207] <= 8'b10000001;  Signal[2][207] <= 8'b00000000; 
 Signal[0][208] <= 8'b00011100;  Signal[1][208] <= 8'b10000001;  Signal[2][208] <= 8'b00000000; 
 Signal[0][209] <= 8'b00011101;  Signal[1][209] <= 8'b10000010;  Signal[2][209] <= 8'b00000000; 
 Signal[0][210] <= 8'b00011101;  Signal[1][210] <= 8'b10000010;  Signal[2][210] <= 8'b00000000; 
 Signal[0][211] <= 8'b00011110;  Signal[1][211] <= 8'b10000010;  Signal[2][211] <= 8'b00000000; 
 Signal[0][212] <= 8'b00011110;  Signal[1][212] <= 8'b10000010;  Signal[2][212] <= 8'b00000000; 
 Signal[0][213] <= 8'b00011111;  Signal[1][213] <= 8'b10000011;  Signal[2][213] <= 8'b00000000; 
 Signal[0][214] <= 8'b00100000;  Signal[1][214] <= 8'b10000011;  Signal[2][214] <= 8'b00000000; 
 Signal[0][215] <= 8'b00100000;  Signal[1][215] <= 8'b10000011;  Signal[2][215] <= 8'b00000000; 
 Signal[0][216] <= 8'b00100001;  Signal[1][216] <= 8'b10000011;  Signal[2][216] <= 8'b00000000; 
 Signal[0][217] <= 8'b00100010;  Signal[1][217] <= 8'b10000100;  Signal[2][217] <= 8'b00000000; 
 Signal[0][218] <= 8'b00100010;  Signal[1][218] <= 8'b10000100;  Signal[2][218] <= 8'b00000000; 
 Signal[0][219] <= 8'b00100011;  Signal[1][219] <= 8'b10000100;  Signal[2][219] <= 8'b00000000; 
 Signal[0][220] <= 8'b00100100;  Signal[1][220] <= 8'b10000100;  Signal[2][220] <= 8'b00000000; 
 Signal[0][221] <= 8'b00100101;  Signal[1][221] <= 8'b10000100;  Signal[2][221] <= 8'b00000000; 
 Signal[0][222] <= 8'b00100101;  Signal[1][222] <= 8'b10000101;  Signal[2][222] <= 8'b00000000; 
 Signal[0][223] <= 8'b00100110;  Signal[1][223] <= 8'b10000101;  Signal[2][223] <= 8'b00000000; 
 Signal[0][224] <= 8'b00100111;  Signal[1][224] <= 8'b10000101;  Signal[2][224] <= 8'b00000000; 
 Signal[0][225] <= 8'b00101000;  Signal[1][225] <= 8'b10000101;  Signal[2][225] <= 8'b00000000; 
 Signal[0][226] <= 8'b00101001;  Signal[1][226] <= 8'b10000101;  Signal[2][226] <= 8'b00000000; 
 Signal[0][227] <= 8'b00101010;  Signal[1][227] <= 8'b10000110;  Signal[2][227] <= 8'b00000000; 
 Signal[0][228] <= 8'b00101011;  Signal[1][228] <= 8'b10000110;  Signal[2][228] <= 8'b00000000; 
 Signal[0][229] <= 8'b00101100;  Signal[1][229] <= 8'b10000110;  Signal[2][229] <= 8'b00000000; 
 Signal[0][230] <= 8'b00101101;  Signal[1][230] <= 8'b10000110;  Signal[2][230] <= 8'b00000000; 
 Signal[0][231] <= 8'b00101110;  Signal[1][231] <= 8'b10000110;  Signal[2][231] <= 8'b00000000; 
 Signal[0][232] <= 8'b00101111;  Signal[1][232] <= 8'b10000110;  Signal[2][232] <= 8'b00000000; 
 Signal[0][233] <= 8'b00110000;  Signal[1][233] <= 8'b10000111;  Signal[2][233] <= 8'b00000000; 
 Signal[0][234] <= 8'b00110001;  Signal[1][234] <= 8'b10000111;  Signal[2][234] <= 8'b00000000; 
 Signal[0][235] <= 8'b00110010;  Signal[1][235] <= 8'b10000111;  Signal[2][235] <= 8'b00000000; 
 Signal[0][236] <= 8'b00110011;  Signal[1][236] <= 8'b10000111;  Signal[2][236] <= 8'b00000000; 
 Signal[0][237] <= 8'b00110100;  Signal[1][237] <= 8'b10000111;  Signal[2][237] <= 8'b00000000; 
 Signal[0][238] <= 8'b00110101;  Signal[1][238] <= 8'b10000111;  Signal[2][238] <= 8'b00000000; 
 Signal[0][239] <= 8'b00110110;  Signal[1][239] <= 8'b10000111;  Signal[2][239] <= 8'b00000000; 
 Signal[0][240] <= 8'b00110111;  Signal[1][240] <= 8'b10001000;  Signal[2][240] <= 8'b00000000; 
 Signal[0][241] <= 8'b00111001;  Signal[1][241] <= 8'b10001000;  Signal[2][241] <= 8'b00000000; 
 Signal[0][242] <= 8'b00111010;  Signal[1][242] <= 8'b10001000;  Signal[2][242] <= 8'b00000000; 
 Signal[0][243] <= 8'b00111011;  Signal[1][243] <= 8'b10001000;  Signal[2][243] <= 8'b00000000; 
 Signal[0][244] <= 8'b00111100;  Signal[1][244] <= 8'b10001000;  Signal[2][244] <= 8'b00000000; 
 Signal[0][245] <= 8'b00111101;  Signal[1][245] <= 8'b10001000;  Signal[2][245] <= 8'b00000000; 
 Signal[0][246] <= 8'b00111110;  Signal[1][246] <= 8'b10001000;  Signal[2][246] <= 8'b00000000; 
 Signal[0][247] <= 8'b01000000;  Signal[1][247] <= 8'b10001001;  Signal[2][247] <= 8'b00000000; 
 Signal[0][248] <= 8'b01000001;  Signal[1][248] <= 8'b10001001;  Signal[2][248] <= 8'b00000000; 
 Signal[0][249] <= 8'b01000010;  Signal[1][249] <= 8'b10001001;  Signal[2][249] <= 8'b00000000; 
 Signal[0][250] <= 8'b01000011;  Signal[1][250] <= 8'b10001001;  Signal[2][250] <= 8'b00000000; 
 Signal[0][251] <= 8'b01000100;  Signal[1][251] <= 8'b10001001;  Signal[2][251] <= 8'b00000000; 
 Signal[0][252] <= 8'b01000110;  Signal[1][252] <= 8'b10001001;  Signal[2][252] <= 8'b00000000; 
 Signal[0][253] <= 8'b01000111;  Signal[1][253] <= 8'b10001001;  Signal[2][253] <= 8'b00000000; 
 Signal[0][254] <= 8'b01001000;  Signal[1][254] <= 8'b10001001;  Signal[2][254] <= 8'b00000000; 
 Signal[0][255] <= 8'b01001001;  Signal[1][255] <= 8'b10001010;  Signal[2][255] <= 8'b00000000; 
 
end  
  


  
endmodule